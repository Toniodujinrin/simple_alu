`ifndef INT_CONVERTER_TEST_SV
`define INT_CONVERTER_TEST_SV 


`ifndef DATA_WIDTH
`define DATA_WIDTH 16
`endif 

module int_converter_testbench; 
    int_converter_interface int_inf(); 
    test tst(int_inf); 
    int_converter DUT(
        .x(int_inf.x), 
        .r(int_inf.r), 
        .negative(int_inf.negative), 
        .cout(int_inf.cout), 
        .overflow(int_inf.overflow), 
        .zero(int_inf.zero)
  );


    initial begin
        $dumpfile("int_converter_test.vcd");
        $dumpvars; 
    end

    initial begin
        #100000;
        $finish;
    end

endmodule:int_converter_testbench


interface int_converter_interface; 
    shortint x;
    bit  [`DATA_WIDTH-1:0] r;
    logic negative; 
    logic zero; 
    logic overflow; 
    logic cout;
endinterface 

class float16;
    bit [9:0] mantissa; 
    bit [4:0] exponent; 
    bit sign;

    function new(bit [15:0] float_val); 
        mantissa = float_val[9:0]; 
        exponent = float_val[14:10]; 
        sign     = float_val[15]; 
    endfunction : new

    function real convert_to_real(); 
        bit implicit_leading_one;
        int real_exponent;
        real frac, result;

        // Special cases
        if (exponent == 5'b0 && mantissa == 10'b0) begin
            return sign ? -0.0 : 0.0;
        end else if (exponent == 5'b11111 && mantissa == 10'b0) begin
            return sign ? -1.0/0.0 : 1.0/0.0; // ±inf
        end else if (exponent == 5'b11111 && mantissa != 10'b0) begin
            return 0.0/0.0; // NaN
        end

        // Normal/denormal
        if (exponent == 0) begin
            real_exponent = -14; // denormal exponent
            implicit_leading_one = 0;
        end else begin
            real_exponent = exponent - 15; // re-bias
            implicit_leading_one = 1;
        end

        // Fraction = implicit + mantissa/1024.0
        frac = implicit_leading_one + (mantissa / 1024.0);

        // Final result
        result = (sign ? -1.0 : 1.0) * (2.0 ** real_exponent) * frac;
        return result;
    endfunction : convert_to_real
endclass : float16



class transaction; 
    rand shortint  x;
    bit  [`DATA_WIDTH-1:0] r; 
    logic negative; 
    logic zero; 
    logic overflow; 
    logic cout;



    function void display();
        float16 r_float = new(r);
        real r_real = r_float.convert_to_real();
      $display("x = %0d, r = %0d, r_raw = %0b  overflow = %0b, negative = %0b, zero = %0b, cout = %0b", x, r_real,r, overflow, negative, zero, cout);
    endfunction:display

endclass: transaction 


class generator; 
    mailbox gen_drv; 
    int samples;
    transaction int_conv_transaction;  

    function new(mailbox gen_drv, int samples); 
        this.gen_drv = gen_drv; 
        this.samples = samples; 
    endfunction: new

    task run(); 
        repeat(samples)
            begin
                int_conv_transaction = new(); 
                assert(int_conv_transaction.randomize()); 
                gen_drv.put(int_conv_transaction); 
            end
    endtask 

endclass:generator


class driver; 
    mailbox gen_drv; 
    int samples; 
    virtual int_converter_interface int_conv_inf; 


  function new(mailbox gen_drv, int samples, virtual int_converter_interface int_conv_inf);
        this.samples = samples; 
        this.gen_drv = gen_drv;
        this.int_conv_inf = int_conv_inf; 
    endfunction:new

    task run();
        repeat(samples)
        begin
          	transaction int_conv_transaction; 
            gen_drv.get(int_conv_transaction); 
            int_conv_inf.x = int_conv_transaction.x; 
            #10; //wait 10 for DUT to process outputs  
        end
    endtask:run

endclass: driver 


class monitor; 
    mailbox mon_sb; 
    int samples; 
    virtual int_converter_interface int_conv_inf; 


    function new(virtual int_converter_interface int_conv_inf, int samples, mailbox mon_sb); 
        this.int_conv_inf = int_conv_inf; 
        this.samples = samples; 
        this.mon_sb = mon_sb; 
    endfunction:new

    task run(); 
        repeat(samples)
        begin
            transaction int_conv_transaction;
            int_conv_transaction = new(); 
            #11; 
            int_conv_transaction.x = int_conv_inf.x; 
            int_conv_transaction.r = int_conv_inf.r; 
            int_conv_transaction.negative = int_conv_inf.negative; 
            int_conv_transaction.zero = int_conv_inf.zero; 
            int_conv_transaction.overflow = int_conv_inf.overflow; 
            int_conv_transaction.cout = int_conv_inf.cout; 
            mon_sb.put(int_conv_transaction); 

        end
    endtask:run

endclass: monitor 


class scoreboard; 
    mailbox mon_sb;
    int samples;
    transaction int_conv_transaction;

    // DUT output
    shortint signed_x; 
    bit [`DATA_WIDTH-1:0] r;
    float16 r_float;
    real r_real; 
    bit overflow, negative, zero, cout;

    // Expected
    shortint expected_x; 
    real expected_r; 
    bit expected_overflow, expected_negative, expected_zero, expected_cout;

    function new(mailbox mon_sb, int samples); 
        this.mon_sb = mon_sb; 
        this.samples = samples; 
    endfunction : new

    task run(); 
        repeat(samples) begin
            mon_sb.get(int_conv_transaction); 

            // DUT output
            signed_x = int_conv_transaction.x;
            r        = int_conv_transaction.r;
            r_float  = new(r);
            r_real   = r_float.convert_to_real();
            overflow = int_conv_transaction.overflow;
            negative = int_conv_transaction.negative;
            zero     = int_conv_transaction.zero;
            cout     = int_conv_transaction.cout;

            // Golden model
            expected_x        = signed_x;
            expected_r        = expected_x; // direct cast to real
            expected_negative = (expected_r < 0);
            expected_zero     = (expected_r == 0);
            expected_overflow = 1'b0; // TODO: implement overflow modeling if needed
            expected_cout     = 1'b0;

            int_conv_transaction.display();

            // Compare results
          if ((expected_r - r_real > 8)|| (expected_r - r_real < -8)) //use an accuracy of +-8 for float comparison
                $error("Int→Float result mismatch: DUT r = %0f, expected r = %0f", r_real, expected_r);
            if (expected_negative !== negative)
                $error("Int→Float negative flag mismatch: DUT negative = %0b, expected = %0b", negative, expected_negative);
            if (expected_zero !== zero) 
                $error("Int→Float zero flag mismatch: DUT zero = %0b, expected = %0b", zero, expected_zero);
            if (expected_overflow !== overflow)
                $error("Int→Float overflow flag mismatch: DUT overflow = %0b, expected = %0b", overflow, expected_overflow);
            if (expected_cout !== cout) 
                $error("Int→Float cout flag mismatch: DUT cout = %0b, expected = %0b", cout, expected_cout);
        end
    endtask : run
endclass : scoreboard


class environment; 
    mailbox gen_drv;
    mailbox mon_sb; 
    int samples; 

    generator gen; 
    driver drv; 
    monitor mon; 
    scoreboard sb; 

    virtual int_converter_interface int_conv_inf;

    function new(virtual int_converter_interface int_conv_inf, int samples); 
        this.int_conv_inf = int_conv_inf; 
        this.samples = samples; 

        gen_drv = new(); 
        mon_sb = new(); 

        gen = new(gen_drv, samples); 
        drv = new(gen_drv, samples, int_conv_inf); 
        mon = new(int_conv_inf, samples, mon_sb); 
        sb = new(mon_sb, samples); 
    endfunction:new

    task run(); 
        fork
            gen.run();
            drv.run();
            mon.run();
            sb.run();
        join
    endtask:run

endclass:environment


program test (int_converter_interface int_conv_inf); 
    int samples = 1000;
    environment env; 
   

    initial begin
        env = new(int_conv_inf, samples); 
        env.run();
    end

endprogram:test


`endif //MULTIPLIER_TEST_SV