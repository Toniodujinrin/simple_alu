module shift(x,y,shift_count,mode, negative, zero, cout, overflow ); 
	parameter WIDTH = 16;
   function integer clogb2;
		input [31:0] value;
		integer 	i;
		begin
			clogb2 = 0;
			for(i = 0; 2**i < value; i = i + 1)
				clogb2 = i + 1;
		end
	endfunction	
	parameter SHIFT_WIDTH = clogb2(WIDTH); 
	input [WIDTH-1:0] x; 
	output [WIDTH-1:0] y; 
	input [SHIFT_WIDTH-1:0] shift_count; 
	input [2:0] mode; 
	//modes////////
	//LSL = 3'b000
	//LSR = 3'b001 
	//ASR = 3'b010 
	//ASL = 3'b011 
	//ROR = 3'b100
	///////////////
	
	wire [WIDTH-1:0] stage_shift [0:SHIFT_WIDTH-1];
	wire [WIDTH-1:0] zero_input = 0;
	wire [WIDTH-1:0] sign_bit_input = {(WIDTH){x[WIDTH-1]}}; 
   
	
	genvar i; 
	generate 
	for(i=0; i < SHIFT_WIDTH; i = i+1)
		begin:BARREL_SHIFT 
			if(i == 0)
					chained_mux#(.WIDTH(WIDTH)) N_MUX(
									 .x(x),
									 .y(
									 mode==3'b100 ? {x[(1 << i)-1:0],x[WIDTH-1:(1 << i)]}: //ROR 
									 mode==3'b001 ? {zero_input[(1 << i)-1:0],x[WIDTH-1:(1 << i)]}:       //LSR
									 mode==3'b010 ? {sign_bit_input[(1 << i)-1:0],x[WIDTH-1:(1 << i)]}:   //ASR
									 mode==3'b000 ? {x[(1 << i)-1:0],zero_input[WIDTH-1:(1 << i)]}: //LSL
									 {x[(1 << i)-1:0],zero_input[WIDTH-1:(1 << i)]} //ASL
									 ), 
									 .s(shift_count[i]),
									 .out(stage_shift[i])); 
			else 
					chained_mux#(.WIDTH(WIDTH)) N_MUX(
									 .x(stage_shift[i-1]),
									 .y(
									 mode==3'b100 ? {stage_shift[i-1][(1 << i)-1:0],stage_shift[i-1][WIDTH-1:(1 << i)]}: //ROR 
									 mode==3'b001 ? {zero_input[(1 << i)-1:0],stage_shift[i-1][WIDTH-1:(1 << i)]}:       //LSR
									 mode==3'b010 ? {sign_bit_input[(1 << i)-1:0],stage_shift[i-1][WIDTH-1:(1 << i)]}:   //ASR
									 mode==3'b000 ? {stage_shift[i-1][(1 << i)-1:0],zero_input[WIDTH-1:(1 << i)]}: //LSL
									 {stage_shift[i-1][(1 << i)-1:0],zero_input[WIDTH-1:(1 << i)]} //ASL
									 ), 
									 .s(shift_count[i]), .out(stage_shift[i])); 
		end 
	endgenerate
	assign y = stage_shift[SHIFT_WIDTH-1]; 
	assign negative = y[WIDTH-1]; 
	assign zero = ~|y; 
	assign cout = 0; 
	assign overflow: (mode == 3'b000) || (mode == 3'b011) && 
	(x[WIDTH-1] ^ Y[WIDTH-1]); 
endmodule 


